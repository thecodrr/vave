module wav

//TODO