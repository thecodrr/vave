module vave

//TODO